module download

pub fn download_song_url(url string) !string {
	return url
}

pub fn download_song_query(query string) !string {
	return query
}

pub fn download_playlist_url(url string) ![]string {
	return [url]
}
